// Адаптер для подключения к мантии Caravel
module user_project_wrapper (
    input  clk,          // Тактовая частота от мантии (10 МГц)
    input  rst_n,        // Сброс от мантии
    
    // Внешние выводы кристалла (ограничено 8 пинами)
    inout  [7:0] io_in,   // Bidirectional пины
    output [7:0] io_out,  // Выходы
    output [7:0] io_oeb   // Направление: 1 = выход, 0 = вход
);

    // Экземпляр вашего счётчика
    counter uut (
        .clk(clk),
        .rst_n(rst_n),
        .count(io_out[3:0])  // Выводим 4 бита на пины 0-3
    );
    
    // Настройка направления пинов:
    // Пины 0-3 = выходы (счётчик), пины 4-7 = входы (не используются)
    assign io_oeb = 8'b11110000;
    
    // Подтягиваем неиспользуемые выходы к 0
    assign io_out[7:4] = 4'b0000;

endmodule
